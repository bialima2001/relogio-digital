library IEEE;
use IEEE.std_logic_1164.ALL;

entity Clock is
	port(clk: in std_logic;
		a0,a1,a2,a3 : out std_logic_vector(3 downto 0)
	);
end;

architecture arq of Clock is
	
	component bcd_7seg_decoder is
		port (
			BCD	: in std_logic_vector(3 downto 0);
			HEX 	: out std_logic_vector(6 downto 0)
		);
	end component;
	
	component contador is
		port(
			bcd	: out std_logic_vector(3 downto 0);
			clk	: in std_logic;
			reset	: in std_logic
		);
	end component;
	
	 
	signal ac0,ac1,ac2,ac3 : std_logic_vector(3 downto 0);
	signal reset0,reset1,reset2,reset3,aux : std_logic;
	
	
begin

a0 <= ac0;
a1 <= ac1;
a2 <= ac2;
a3 <= ac3;

		
counter0 : contador
	port map(ac0,clk,reset0);
	
reset0 <= '1' when ac0 = x"A" else '0';
	
counter1 : contador
	port map(ac1,reset0,reset1);
	
reset1 <= '1' when ac1 = x"6" else '0';
	
counter2 : contador
	port map(
		ac2,
		reset1,
		reset2
	);

reset2 <=
	'1' when ac2 = x"A" else
	'1' when ac3 = x"2" and ac2 = x"4" else
	'0';
	
aux <= '1' when ac2 = x"A" else '0';

counter3 : contador
	port map(ac3,aux,reset3);
	

reset3 <=
	'1' when ac3 = x"2" and ac2 = x"4" else
	'0';

end;
